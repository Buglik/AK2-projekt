VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO full_adder
   CLASS BLOCK ;
   FOREIGN full_adder ;
   ORIGIN 2.6000 -0.0000 ;
   SIZE 38.7000 BY 13.1000 ;
   PIN vdd
      PORT
         LAYER metal1 ;
	    RECT 0.6000 0.8000 1.0000 3.1000 ;
	    RECT 2.2000 0.8000 2.6000 4.9000 ;
	    RECT 5.4000 0.8000 5.8000 5.1000 ;
	    RECT 6.2000 0.8000 6.6000 3.1000 ;
	    RECT 7.8000 0.8000 8.2000 3.1000 ;
	    RECT 11.5000 0.8000 11.9000 5.1000 ;
	    RECT 14.2000 0.8000 14.6000 2.9000 ;
	    RECT 15.8000 0.8000 16.2000 3.1000 ;
	    RECT 16.9000 0.8000 17.3000 3.1000 ;
	    RECT 19.0000 0.8000 19.4000 5.1000 ;
	    RECT 20.6000 0.8000 21.0000 3.1000 ;
	    RECT 21.4000 0.8000 21.8000 5.1000 ;
	    RECT 23.5000 0.8000 23.9000 3.1000 ;
	    RECT 26.2000 0.8000 26.6000 3.1000 ;
	    RECT 27.8000 0.8000 28.2000 3.1000 ;
	    RECT 29.4000 0.8000 29.8000 4.5000 ;
	    RECT 31.8000 0.8000 32.2000 4.5000 ;
	    RECT 0.2000 0.2000 33.4000 0.8000 ;
         LAYER metal2 ;
	    RECT 8.0000 0.3000 9.6000 0.7000 ;
         LAYER metal3 ;
	    RECT 8.0000 0.3000 9.6000 0.7000 ;
         LAYER metal4 ;
	    RECT 8.0000 0.3000 9.6000 0.7000 ;
         LAYER metal5 ;
	    RECT 8.0000 0.7000 8.6000 0.8000 ;
	    RECT 9.0000 0.7000 9.6000 0.8000 ;
	    RECT 8.0000 0.2000 9.6000 0.7000 ;
         LAYER metal6 ;
	    RECT 8.0000 0.0000 9.6000 13.0000 ;
      END
   END vdd
   PIN gnd
      PORT
         LAYER metal1 ;
	    RECT 0.2000 10.2000 33.4000 10.8000 ;
	    RECT 1.9000 8.0000 2.3000 10.2000 ;
	    RECT 3.8000 8.9000 4.2000 10.2000 ;
	    RECT 5.4000 8.9000 5.8000 10.2000 ;
	    RECT 6.2000 7.9000 6.6000 10.2000 ;
	    RECT 10.2000 8.9000 10.6000 10.2000 ;
	    RECT 11.8000 8.1000 12.2000 10.2000 ;
	    RECT 15.8000 6.9000 16.2000 10.2000 ;
	    RECT 18.2000 8.3000 18.6000 10.2000 ;
	    RECT 20.6000 8.9000 21.0000 10.2000 ;
	    RECT 22.2000 8.3000 22.6000 10.2000 ;
	    RECT 26.2000 7.9000 26.6000 10.2000 ;
	    RECT 29.4000 7.9000 29.8000 10.2000 ;
	    RECT 31.8000 7.9000 32.2000 10.2000 ;
         LAYER metal2 ;
	    RECT 24.0000 10.3000 25.6000 10.7000 ;
         LAYER metal3 ;
	    RECT 24.0000 10.3000 25.6000 10.7000 ;
         LAYER metal4 ;
	    RECT 24.0000 10.3000 25.6000 10.7000 ;
         LAYER metal5 ;
	    RECT 24.0000 10.7000 24.6000 10.8000 ;
	    RECT 25.0000 10.7000 25.6000 10.8000 ;
	    RECT 24.0000 10.2000 25.6000 10.7000 ;
         LAYER metal6 ;
	    RECT 24.0000 0.0000 25.6000 13.0000 ;
      END
   END gnd
   PIN i_x
      PORT
         LAYER metal1 ;
	    RECT 7.8000 7.1000 8.2000 7.2000 ;
	    RECT 11.0000 7.1000 11.5000 7.2000 ;
	    RECT 1.6000 6.9000 2.0000 7.0000 ;
	    RECT 1.5000 6.6000 2.0000 6.9000 ;
	    RECT 7.8000 6.8000 11.5000 7.1000 ;
	    RECT 1.5000 6.2000 1.8000 6.6000 ;
	    RECT 11.2000 6.4000 11.6000 6.8000 ;
	    RECT 1.4000 5.8000 1.8000 6.2000 ;
	    RECT 3.8000 5.4000 4.2000 6.2000 ;
	    RECT 7.8000 4.4000 8.2000 5.2000 ;
         LAYER metal2 ;
	    RECT 1.4000 6.8000 1.8000 7.2000 ;
	    RECT 3.8000 6.8000 4.2000 7.2000 ;
	    RECT 7.8000 6.8000 8.2000 7.2000 ;
	    RECT 1.4000 6.2000 1.7000 6.8000 ;
	    RECT 3.8000 6.2000 4.1000 6.8000 ;
	    RECT 7.8000 6.2000 8.1000 6.8000 ;
	    RECT 1.4000 5.8000 1.8000 6.2000 ;
	    RECT 3.8000 5.8000 4.2000 6.2000 ;
	    RECT 7.8000 5.8000 8.2000 6.2000 ;
	    RECT 7.8000 5.2000 8.1000 5.8000 ;
	    RECT 7.8000 4.8000 8.2000 5.2000 ;
         LAYER metal3 ;
	    RECT 1.4000 6.8000 1.8000 7.2000 ;
	    RECT 3.8000 6.8000 4.2000 7.2000 ;
	    RECT 1.4000 6.1000 1.7000 6.8000 ;
	    RECT 3.8000 6.1000 4.1000 6.8000 ;
	    RECT 7.8000 6.1000 8.2000 6.2000 ;
	    RECT -2.6000 5.8000 8.2000 6.1000 ;
      END
   END i_x
   PIN i_y
      PORT
         LAYER metal1 ;
	    RECT 5.4000 7.8000 5.8000 8.6000 ;
	    RECT 8.6000 8.1000 9.0000 8.2000 ;
	    RECT 10.2000 8.1000 10.6000 8.6000 ;
	    RECT 8.6000 7.8000 10.6000 8.1000 ;
	    RECT 0.6000 6.4000 1.0000 7.2000 ;
	    RECT 5.4000 7.1000 5.7000 7.8000 ;
	    RECT 6.2000 7.1000 6.6000 7.6000 ;
	    RECT 5.4000 6.8000 6.6000 7.1000 ;
         LAYER metal2 ;
	    RECT 0.6000 7.8000 1.0000 8.2000 ;
	    RECT 6.2000 7.8000 6.6000 8.2000 ;
	    RECT 8.6000 7.8000 9.0000 8.2000 ;
	    RECT 0.6000 7.2000 0.9000 7.8000 ;
	    RECT 6.2000 7.2000 6.5000 7.8000 ;
	    RECT 8.6000 7.2000 8.9000 7.8000 ;
	    RECT 0.6000 6.8000 1.0000 7.2000 ;
	    RECT 6.2000 7.1000 6.6000 7.2000 ;
	    RECT 7.0000 7.1000 7.4000 7.2000 ;
	    RECT 6.2000 6.8000 7.4000 7.1000 ;
	    RECT 8.6000 6.8000 9.0000 7.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 8.1000 1.0000 8.2000 ;
	    RECT 6.2000 8.1000 6.6000 8.2000 ;
	    RECT -2.6000 7.8000 6.6000 8.1000 ;
	    RECT 7.0000 7.1000 7.4000 7.2000 ;
	    RECT 8.6000 7.1000 9.0000 7.2000 ;
	    RECT 7.0000 6.8000 9.0000 7.1000 ;
      END
   END i_y
   PIN i_carry
      PORT
         LAYER metal1 ;
	    RECT 20.6000 7.8000 21.0000 8.6000 ;
	    RECT 23.8000 5.1000 24.2000 5.2000 ;
	    RECT 23.5000 4.8000 24.2000 5.1000 ;
	    RECT 23.5000 4.2000 23.8000 4.8000 ;
	    RECT 23.4000 3.8000 23.8000 4.2000 ;
         LAYER metal2 ;
	    RECT 20.6000 9.2000 20.9000 13.1000 ;
	    RECT 20.6000 8.8000 21.0000 9.2000 ;
	    RECT 23.8000 8.8000 24.2000 9.2000 ;
	    RECT 20.6000 8.2000 20.9000 8.8000 ;
	    RECT 20.6000 7.8000 21.0000 8.2000 ;
	    RECT 23.8000 5.2000 24.1000 8.8000 ;
	    RECT 23.8000 4.8000 24.2000 5.2000 ;
         LAYER metal3 ;
	    RECT 20.6000 9.1000 21.0000 9.2000 ;
	    RECT 23.8000 9.1000 24.2000 9.2000 ;
	    RECT 20.6000 8.8000 24.2000 9.1000 ;
      END
   END i_carry
   PIN o_sum
      PORT
         LAYER metal1 ;
	    RECT 30.2000 6.2000 30.6000 9.9000 ;
	    RECT 30.3000 5.1000 30.6000 6.2000 ;
	    RECT 30.2000 1.1000 30.6000 5.1000 ;
         LAYER metal2 ;
	    RECT 30.2000 8.8000 30.6000 9.2000 ;
	    RECT 30.2000 8.2000 30.5000 8.8000 ;
	    RECT 30.2000 7.8000 30.6000 8.2000 ;
         LAYER metal3 ;
	    RECT 30.2000 8.8000 30.6000 9.2000 ;
	    RECT 30.2000 8.1000 30.5000 8.8000 ;
	    RECT 30.2000 7.8000 36.1000 8.1000 ;
      END
   END o_sum
   PIN o_carry
      PORT
         LAYER metal1 ;
	    RECT 32.6000 6.2000 33.0000 9.9000 ;
	    RECT 32.7000 5.1000 33.0000 6.2000 ;
	    RECT 32.6000 1.1000 33.0000 5.1000 ;
         LAYER metal2 ;
	    RECT 32.6000 6.8000 33.0000 7.2000 ;
	    RECT 32.6000 6.2000 32.9000 6.8000 ;
	    RECT 32.6000 5.8000 33.0000 6.2000 ;
         LAYER metal3 ;
	    RECT 32.6000 6.1000 33.0000 6.2000 ;
	    RECT 32.6000 5.8000 36.1000 6.1000 ;
      END
   END o_carry
   OBS
         LAYER metal1 ;
	    RECT 0.6000 7.9000 1.0000 9.9000 ;
	    RECT 2.7000 8.4000 3.1000 9.9000 ;
	    RECT 4.6000 8.9000 5.0000 9.9000 ;
	    RECT 2.7000 7.9000 3.4000 8.4000 ;
	    RECT 0.7000 7.8000 1.0000 7.9000 ;
	    RECT 0.7000 7.6000 1.6000 7.8000 ;
	    RECT 0.7000 7.5000 2.8000 7.6000 ;
	    RECT 1.3000 7.3000 2.8000 7.5000 ;
	    RECT 2.4000 7.2000 2.8000 7.3000 ;
	    RECT 2.4000 5.5000 2.7000 7.2000 ;
	    RECT 3.1000 6.2000 3.4000 7.9000 ;
	    RECT 3.0000 5.8000 3.4000 6.2000 ;
	    RECT 1.5000 5.2000 2.7000 5.5000 ;
	    RECT 1.5000 3.1000 1.8000 5.2000 ;
	    RECT 3.1000 5.1000 3.4000 5.8000 ;
	    RECT 4.6000 7.2000 4.9000 8.9000 ;
	    RECT 7.5000 8.2000 7.9000 9.9000 ;
	    RECT 11.0000 8.9000 11.4000 9.9000 ;
	    RECT 7.0000 7.9000 7.9000 8.2000 ;
	    RECT 4.6000 6.8000 5.0000 7.2000 ;
	    RECT 4.6000 5.2000 4.9000 6.8000 ;
	    RECT 7.0000 6.1000 7.4000 7.9000 ;
	    RECT 11.1000 7.8000 11.4000 8.9000 ;
	    RECT 12.6000 7.9000 13.0000 9.9000 ;
	    RECT 11.1000 7.5000 12.3000 7.8000 ;
	    RECT 8.6000 6.1000 9.0000 6.2000 ;
	    RECT 7.0000 5.8000 9.0000 6.1000 ;
	    RECT 12.0000 6.0000 12.3000 7.5000 ;
	    RECT 12.7000 6.2000 13.0000 7.9000 ;
	    RECT 14.0000 7.1000 14.4000 9.9000 ;
	    RECT 16.6000 7.9000 17.0000 9.9000 ;
	    RECT 17.4000 8.0000 17.8000 9.9000 ;
	    RECT 19.0000 8.0000 19.4000 9.9000 ;
	    RECT 17.4000 7.9000 19.4000 8.0000 ;
	    RECT 16.7000 7.2000 17.0000 7.9000 ;
	    RECT 17.5000 7.7000 19.3000 7.9000 ;
	    RECT 18.6000 7.2000 19.0000 7.4000 ;
	    RECT 4.6000 5.1000 5.0000 5.2000 ;
	    RECT 1.4000 1.1000 1.8000 3.1000 ;
	    RECT 3.0000 1.1000 3.4000 5.1000 ;
	    RECT 4.1000 4.7000 5.0000 5.1000 ;
	    RECT 4.1000 1.1000 4.5000 4.7000 ;
	    RECT 7.0000 1.1000 7.4000 5.8000 ;
	    RECT 11.9000 5.7000 12.3000 6.0000 ;
	    RECT 12.6000 5.8000 13.0000 6.2000 ;
	    RECT 10.2000 5.6000 12.3000 5.7000 ;
	    RECT 10.2000 5.4000 12.2000 5.6000 ;
	    RECT 10.2000 1.1000 10.6000 5.4000 ;
	    RECT 12.7000 5.1000 13.0000 5.8000 ;
	    RECT 13.5000 6.9000 14.4000 7.1000 ;
	    RECT 13.5000 6.8000 14.3000 6.9000 ;
	    RECT 16.6000 6.8000 17.9000 7.2000 ;
	    RECT 18.6000 6.9000 19.4000 7.2000 ;
	    RECT 19.0000 6.8000 19.4000 6.9000 ;
	    RECT 13.5000 5.2000 13.8000 6.8000 ;
	    RECT 14.6000 5.8000 15.4000 6.2000 ;
	    RECT 12.3000 4.8000 13.0000 5.1000 ;
	    RECT 13.4000 4.8000 13.8000 5.2000 ;
	    RECT 15.8000 4.8000 16.2000 6.2000 ;
	    RECT 16.6000 5.1000 17.0000 5.2000 ;
	    RECT 17.6000 5.1000 17.9000 6.8000 ;
	    RECT 18.2000 6.1000 18.6000 6.6000 ;
	    RECT 19.8000 6.1000 20.2000 9.9000 ;
	    RECT 21.4000 8.0000 21.8000 9.9000 ;
	    RECT 23.0000 8.0000 23.4000 9.9000 ;
	    RECT 21.4000 7.9000 23.4000 8.0000 ;
	    RECT 23.8000 7.9000 24.2000 9.9000 ;
	    RECT 27.5000 8.2000 27.9000 9.9000 ;
	    RECT 27.0000 7.9000 27.9000 8.2000 ;
	    RECT 21.5000 7.7000 23.3000 7.9000 ;
	    RECT 21.8000 7.2000 22.2000 7.4000 ;
	    RECT 23.8000 7.2000 24.1000 7.9000 ;
	    RECT 21.4000 6.9000 22.2000 7.2000 ;
	    RECT 22.9000 7.1000 24.2000 7.2000 ;
	    RECT 26.2000 7.1000 26.6000 7.6000 ;
	    RECT 21.4000 6.8000 21.8000 6.9000 ;
	    RECT 22.9000 6.8000 26.6000 7.1000 ;
	    RECT 18.2000 5.8000 20.2000 6.1000 ;
	    RECT 22.2000 5.8000 22.6000 6.6000 ;
	    RECT 16.6000 4.8000 17.3000 5.1000 ;
	    RECT 17.6000 4.8000 18.1000 5.1000 ;
	    RECT 12.3000 4.2000 12.7000 4.8000 ;
	    RECT 12.3000 3.8000 13.0000 4.2000 ;
	    RECT 12.3000 1.1000 12.7000 3.8000 ;
	    RECT 13.5000 3.5000 13.8000 4.8000 ;
	    RECT 14.2000 3.8000 14.6000 4.6000 ;
	    RECT 17.0000 4.2000 17.3000 4.8000 ;
	    RECT 17.0000 3.8000 17.4000 4.2000 ;
	    RECT 13.5000 3.2000 15.3000 3.5000 ;
	    RECT 17.7000 3.2000 18.1000 4.8000 ;
	    RECT 13.5000 3.1000 13.8000 3.2000 ;
	    RECT 13.4000 1.1000 13.8000 3.1000 ;
	    RECT 15.0000 1.1000 15.4000 3.2000 ;
	    RECT 17.7000 2.8000 18.6000 3.2000 ;
	    RECT 17.7000 1.1000 18.1000 2.8000 ;
	    RECT 19.8000 1.1000 20.2000 5.8000 ;
	    RECT 22.9000 5.1000 23.2000 6.8000 ;
	    RECT 22.7000 4.8000 23.2000 5.1000 ;
	    RECT 27.0000 6.1000 27.4000 7.9000 ;
	    RECT 28.6000 7.6000 29.0000 9.9000 ;
	    RECT 31.0000 7.6000 31.4000 9.9000 ;
	    RECT 28.6000 7.3000 29.7000 7.6000 ;
	    RECT 31.0000 7.3000 32.1000 7.6000 ;
	    RECT 28.6000 6.1000 29.0000 6.6000 ;
	    RECT 27.0000 5.8000 29.0000 6.1000 ;
	    RECT 29.4000 5.8000 29.7000 7.3000 ;
	    RECT 31.0000 5.8000 31.4000 6.6000 ;
	    RECT 31.8000 5.8000 32.1000 7.3000 ;
	    RECT 22.7000 1.1000 23.1000 4.8000 ;
	    RECT 27.0000 1.1000 27.4000 5.8000 ;
	    RECT 29.4000 5.4000 30.0000 5.8000 ;
	    RECT 31.8000 5.4000 32.4000 5.8000 ;
	    RECT 27.8000 4.4000 28.2000 5.2000 ;
	    RECT 29.4000 5.1000 29.7000 5.4000 ;
	    RECT 31.8000 5.1000 32.1000 5.4000 ;
	    RECT 28.6000 4.8000 29.7000 5.1000 ;
	    RECT 31.0000 4.8000 32.1000 5.1000 ;
	    RECT 28.6000 1.1000 29.0000 4.8000 ;
	    RECT 31.0000 1.1000 31.4000 4.8000 ;
         LAYER metal2 ;
	    RECT 3.0000 6.8000 3.4000 7.2000 ;
	    RECT 15.8000 6.8000 16.2000 7.2000 ;
	    RECT 18.2000 6.8000 18.6000 7.2000 ;
	    RECT 19.0000 6.8000 19.4000 7.2000 ;
	    RECT 20.6000 7.1000 21.0000 7.2000 ;
	    RECT 21.4000 7.1000 21.8000 7.2000 ;
	    RECT 20.6000 6.8000 21.8000 7.1000 ;
	    RECT 3.0000 6.2000 3.3000 6.8000 ;
	    RECT 15.8000 6.2000 16.1000 6.8000 ;
	    RECT 18.2000 6.2000 18.5000 6.8000 ;
	    RECT 3.0000 5.8000 3.4000 6.2000 ;
	    RECT 8.6000 6.1000 9.0000 6.2000 ;
	    RECT 9.4000 6.1000 9.8000 6.2000 ;
	    RECT 8.6000 5.8000 9.8000 6.1000 ;
	    RECT 14.2000 6.1000 14.6000 6.2000 ;
	    RECT 15.0000 6.1000 15.4000 6.2000 ;
	    RECT 14.2000 5.8000 15.4000 6.1000 ;
	    RECT 15.8000 5.8000 16.2000 6.2000 ;
	    RECT 16.6000 5.8000 17.0000 6.2000 ;
	    RECT 18.2000 5.8000 18.6000 6.2000 ;
	    RECT 16.6000 5.2000 16.9000 5.8000 ;
	    RECT 19.0000 5.2000 19.3000 6.8000 ;
	    RECT 22.2000 5.8000 22.6000 6.2000 ;
	    RECT 31.0000 5.8000 31.4000 6.2000 ;
	    RECT 22.2000 5.2000 22.5000 5.8000 ;
	    RECT 4.6000 4.8000 5.0000 5.2000 ;
	    RECT 16.6000 4.8000 17.0000 5.2000 ;
	    RECT 19.0000 4.8000 19.4000 5.2000 ;
	    RECT 22.2000 4.8000 22.6000 5.2000 ;
	    RECT 27.8000 4.8000 28.2000 5.2000 ;
	    RECT 4.6000 4.2000 4.9000 4.8000 ;
	    RECT 27.8000 4.2000 28.1000 4.8000 ;
	    RECT 4.6000 3.8000 5.0000 4.2000 ;
	    RECT 12.6000 3.8000 13.0000 4.2000 ;
	    RECT 13.4000 4.1000 13.8000 4.2000 ;
	    RECT 14.2000 4.1000 14.6000 4.2000 ;
	    RECT 13.4000 3.8000 14.6000 4.1000 ;
	    RECT 15.0000 3.8000 15.4000 4.2000 ;
	    RECT 27.8000 3.8000 28.2000 4.2000 ;
	    RECT 12.6000 3.2000 12.9000 3.8000 ;
	    RECT 15.0000 3.2000 15.3000 3.8000 ;
	    RECT 31.0000 3.2000 31.3000 5.8000 ;
	    RECT 12.6000 2.8000 13.0000 3.2000 ;
	    RECT 15.0000 2.8000 15.4000 3.2000 ;
	    RECT 18.2000 2.8000 18.6000 3.2000 ;
	    RECT 31.0000 2.8000 31.4000 3.2000 ;
	    RECT 18.2000 2.2000 18.5000 2.8000 ;
	    RECT 18.2000 1.8000 18.6000 2.2000 ;
         LAYER metal3 ;
	    RECT 2.2000 7.1000 2.6000 7.2000 ;
	    RECT 3.0000 7.1000 3.4000 7.2000 ;
	    RECT 2.2000 6.8000 3.4000 7.1000 ;
	    RECT 15.8000 7.1000 16.2000 7.2000 ;
	    RECT 18.2000 7.1000 18.6000 7.2000 ;
	    RECT 15.8000 6.8000 18.6000 7.1000 ;
	    RECT 19.8000 7.1000 20.2000 7.2000 ;
	    RECT 20.6000 7.1000 21.0000 7.2000 ;
	    RECT 19.8000 6.8000 21.0000 7.1000 ;
	    RECT 9.4000 6.1000 9.8000 6.2000 ;
	    RECT 14.2000 6.1000 14.6000 6.2000 ;
	    RECT 16.6000 6.1000 17.0000 6.2000 ;
	    RECT 9.4000 5.8000 17.0000 6.1000 ;
	    RECT 19.0000 5.1000 19.4000 5.2000 ;
	    RECT 22.2000 5.1000 22.6000 5.2000 ;
	    RECT 4.6000 4.8000 22.6000 5.1000 ;
	    RECT 4.6000 4.2000 4.9000 4.8000 ;
	    RECT 4.6000 3.8000 5.0000 4.2000 ;
	    RECT 13.4000 4.1000 13.8000 4.2000 ;
	    RECT 12.6000 3.8000 13.8000 4.1000 ;
	    RECT 15.0000 4.1000 15.4000 4.2000 ;
	    RECT 27.8000 4.1000 28.2000 4.2000 ;
	    RECT 15.0000 3.8000 28.2000 4.1000 ;
	    RECT 12.6000 3.2000 12.9000 3.8000 ;
	    RECT 12.6000 2.8000 13.0000 3.2000 ;
	    RECT 31.0000 3.1000 31.4000 3.2000 ;
	    RECT 18.2000 2.8000 31.4000 3.1000 ;
	    RECT 18.2000 2.2000 18.5000 2.8000 ;
	    RECT 18.2000 1.8000 18.6000 2.2000 ;
         LAYER metal4 ;
	    RECT 2.2000 7.1000 2.6000 7.2000 ;
	    RECT 3.0000 7.1000 3.4000 7.2000 ;
	    RECT 2.2000 6.8000 3.4000 7.1000 ;
	    RECT 19.0000 7.1000 19.4000 7.2000 ;
	    RECT 19.8000 7.1000 20.2000 7.2000 ;
	    RECT 19.0000 6.8000 20.2000 7.1000 ;
         LAYER metal5 ;
	    RECT 3.0000 7.1000 3.4000 7.2000 ;
	    RECT 19.0000 7.1000 19.4000 7.2000 ;
	    RECT 3.0000 6.8000 19.4000 7.1000 ;
   END
END full_adder
