* NGSPICE file created from full_adder.ext - technology: scmos

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

.subckt full_adder vdd gnd i_x i_y i_carry o_sum o_carry
XNAND2X1_2 OAI21X1_1/Y NAND3X1_1/Y gnd BUFX2_2/A vdd NAND2X1
XNOR2X1_1 i_y i_x gnd NOR2X1_1/Y vdd NOR2X1
XOR2X2_1 i_y i_x gnd OR2X2_1/Y vdd OR2X2
XNAND3X1_1 INVX1_1/Y NAND2X1_1/Y OR2X2_1/Y gnd NAND3X1_1/Y vdd NAND3X1
XINVX1_1 i_carry gnd INVX1_1/Y vdd INVX1
XAND2X2_1 i_y i_x gnd AND2X2_1/Y vdd AND2X2
XFILL_0_1_0 gnd vdd FILL
XOAI21X1_1 AND2X2_1/Y NOR2X1_1/Y i_carry gnd OAI21X1_1/Y vdd OAI21X1
XFILL_0_1_1 gnd vdd FILL
XOAI21X1_2 NOR2X1_1/Y INVX1_1/Y NAND2X1_1/Y gnd BUFX2_1/A vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd o_carry vdd BUFX2
XFILL_0_0_0 gnd vdd FILL
XBUFX2_2 BUFX2_2/A gnd o_sum vdd BUFX2
XFILL_0_0_1 gnd vdd FILL
XNAND2X1_1 i_y i_x gnd NAND2X1_1/Y vdd NAND2X1
.ends

