magic
tech scmos
timestamp 1623333969
<< metal1 >>
rect 240 103 242 107
rect 246 103 249 107
rect 253 103 256 107
rect 54 71 57 81
rect 90 78 105 81
rect 54 68 62 71
rect 82 68 113 71
rect 238 68 265 71
rect 70 58 86 61
rect 186 58 201 61
rect 270 58 289 61
rect 158 56 162 58
rect 181 28 182 32
rect 80 3 82 7
rect 86 3 89 7
rect 93 3 96 7
<< m2contact >>
rect 242 103 246 107
rect 249 103 253 107
rect 6 68 10 72
rect 86 78 90 82
rect 206 78 210 82
rect 302 78 306 82
rect 62 68 66 72
rect 78 68 82 72
rect 190 68 194 72
rect 214 68 218 72
rect 326 68 330 72
rect 14 58 18 62
rect 30 58 34 62
rect 38 58 42 62
rect 86 58 90 62
rect 150 58 154 62
rect 158 58 162 62
rect 182 58 186 62
rect 222 58 226 62
rect 310 58 314 62
rect 46 48 50 52
rect 78 48 82 52
rect 166 48 170 52
rect 238 48 242 52
rect 278 48 282 52
rect 126 38 130 42
rect 142 38 146 42
rect 150 28 154 32
rect 182 28 186 32
rect 82 3 86 7
rect 89 3 93 7
<< metal2 >>
rect 206 92 209 131
rect 240 103 242 107
rect 246 103 249 107
rect 253 103 256 107
rect 206 82 209 88
rect 6 72 9 78
rect 62 72 65 78
rect 86 72 89 78
rect 66 68 70 71
rect 210 68 214 71
rect 14 62 17 68
rect 30 62 33 68
rect 38 62 41 68
rect 78 62 81 68
rect 158 62 161 68
rect 182 62 185 68
rect 90 58 94 61
rect 146 58 150 61
rect 78 52 81 58
rect 166 52 169 58
rect 190 52 193 68
rect 222 52 225 58
rect 238 52 241 88
rect 302 82 305 88
rect 326 62 329 68
rect 46 42 49 48
rect 278 42 281 48
rect 138 38 142 41
rect 126 32 129 38
rect 150 32 153 38
rect 310 32 313 58
rect 182 22 185 28
rect 80 3 82 7
rect 86 3 89 7
rect 93 3 96 7
<< m3contact >>
rect 242 103 246 107
rect 249 103 253 107
rect 206 88 210 92
rect 238 88 242 92
rect 302 88 306 92
rect 6 78 10 82
rect 62 78 66 82
rect 14 68 18 72
rect 30 68 34 72
rect 38 68 42 72
rect 70 68 74 72
rect 86 68 90 72
rect 158 68 162 72
rect 182 68 186 72
rect 206 68 210 72
rect 78 58 82 62
rect 94 58 98 62
rect 142 58 146 62
rect 166 58 170 62
rect 326 58 330 62
rect 190 48 194 52
rect 222 48 226 52
rect 46 38 50 42
rect 134 38 138 42
rect 150 38 154 42
rect 278 38 282 42
rect 126 28 130 32
rect 310 28 314 32
rect 182 18 186 22
rect 82 3 86 7
rect 89 3 93 7
<< metal3 >>
rect 240 103 242 107
rect 246 103 249 107
rect 254 103 256 107
rect 210 88 238 91
rect -26 78 6 81
rect 10 78 62 81
rect 302 81 305 88
rect 302 78 361 81
rect 26 68 30 71
rect 74 68 86 71
rect 162 68 182 71
rect 202 68 206 71
rect 14 61 17 68
rect 38 61 41 68
rect -26 58 78 61
rect 98 58 142 61
rect 146 58 166 61
rect 330 58 361 61
rect 46 48 190 51
rect 194 48 222 51
rect 46 42 49 48
rect 126 38 134 41
rect 154 38 278 41
rect 126 32 129 38
rect 182 28 310 31
rect 182 22 185 28
rect 80 3 82 7
rect 86 3 89 7
rect 94 3 96 7
<< m4contact >>
rect 242 103 246 107
rect 250 103 253 107
rect 253 103 254 107
rect 22 68 26 72
rect 198 68 202 72
rect 82 3 86 7
rect 90 3 93 7
rect 93 3 94 7
<< metal4 >>
rect 240 103 242 107
rect 246 103 249 107
rect 254 103 256 107
rect 26 68 30 71
rect 194 68 198 71
rect 80 3 82 7
rect 86 3 89 7
rect 94 3 96 7
<< m5contact >>
rect 242 103 246 107
rect 249 103 250 107
rect 250 103 253 107
rect 30 68 34 72
rect 190 68 194 72
rect 82 3 86 7
rect 89 3 90 7
rect 90 3 93 7
<< metal5 >>
rect 246 103 249 107
rect 246 102 250 103
rect 34 68 190 71
rect 86 3 89 7
rect 86 2 90 3
<< m6contact >>
rect 240 107 246 108
rect 250 107 256 108
rect 240 103 242 107
rect 242 103 246 107
rect 250 103 253 107
rect 253 103 256 107
rect 240 102 246 103
rect 250 102 256 103
rect 80 7 86 8
rect 90 7 96 8
rect 80 3 82 7
rect 82 3 86 7
rect 90 3 93 7
rect 93 3 96 7
rect 80 2 86 3
rect 90 2 96 3
<< metal6 >>
rect 80 8 96 130
rect 86 2 90 8
rect 80 0 96 2
rect 240 108 256 130
rect 246 102 250 108
rect 240 0 256 102
use AND2X2  AND2X2_1
timestamp 1623333969
transform 1 0 4 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_1
timestamp 1623333969
transform -1 0 60 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_1
timestamp 1623333969
transform 1 0 60 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_0_0
timestamp 1623333969
transform 1 0 84 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1623333969
transform 1 0 92 0 -1 105
box -2 -3 10 103
use OR2X2  OR2X2_1
timestamp 1623333969
transform 1 0 100 0 -1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_1
timestamp 1623333969
transform -1 0 164 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_2
timestamp 1623333969
transform -1 0 196 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_1
timestamp 1623333969
transform -1 0 212 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_1
timestamp 1623333969
transform 1 0 212 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_1_0
timestamp 1623333969
transform 1 0 244 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1623333969
transform 1 0 252 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_2
timestamp 1623333969
transform 1 0 260 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_2
timestamp 1623333969
transform 1 0 284 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_1
timestamp 1623333969
transform 1 0 308 0 -1 105
box -2 -3 26 103
<< labels >>
flabel metal6 s 80 0 96 8 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 240 0 256 8 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -24 60 -24 60 7 FreeSans 24 270 0 0 i_x
port 2 nsew
flabel metal3 s -24 80 -24 80 7 FreeSans 24 270 0 0 i_y
port 3 nsew
flabel metal2 s 208 130 208 130 3 FreeSans 24 90 0 0 i_carry
port 4 nsew
flabel metal3 s 360 80 360 80 3 FreeSans 24 270 0 0 o_sum
port 5 nsew
flabel metal3 s 360 60 360 60 3 FreeSans 24 270 0 0 o_carry
port 6 nsew
<< end >>
